----------------------------------------------------------------------------------
-- Company: Nameless2
-- Engineer: Ana María Martínez Gómez, Aitor Alonso Lorenzo, Víctor Adolfo Gallego Alcalá
--
-- Create Date:    16:20:31 02/20/2014 
-- Design Name: 
-- Module Name:    logaritmo - Behavioral 
-- Project Name: Representación gráfica de funciones	
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity logaritmo is
    Port ( valor : in  STD_LOGIC_VECTOR (20 downto 0);
           log : out  STD_LOGIC_VECTOR (20 downto 0);
		   xlogmx : out  STD_LOGIC_VECTOR (20 downto 0));
end logaritmo;

architecture Behavioral of logaritmo is

begin

with valor select
	log 			<=  
"111111111001000100011" when "000000000000000100000",
"111111111010011101000" when "000000000000001000000",
"111111111011010001000" when "000000000000001100000",
"111111111011110101110" when "000000000000010000000",
"111111111100010010011" when "000000000000010100000",
"111111111100101001101" when "000000000000011000000",
"111111111100111101011" when "000000000000011100000",
"111111111101001110100" when "000000000000100000000",
"111111111101011101101" when "000000000000100100000",
"111111111101101011000" when "000000000000101000000",
"111111111101110111010" when "000000000000101100000",
"111111111110000010011" when "000000000000110000000",
"111111111110001100101" when "000000000000110100000",
"111111111110010110001" when "000000000000111000000",
"111111111110011111000" when "000000000000111100000",
"111111111110100111010" when "000000000001000000000",
"111111111110101111000" when "000000000001000100000",
"111111111110110110010" when "000000000001001000000",
"111111111110111101010" when "000000000001001100000",
"111111111111000011110" when "000000000001010000000",
"111111111111001010000" when "000000000001010100000",
"111111111111010000000" when "000000000001011000000",
"111111111111010101101" when "000000000001011100000",
"111111111111011011001" when "000000000001100000000",
"111111111111100000011" when "000000000001100100000",
"111111111111100101011" when "000000000001101000000",
"111111111111101010010" when "000000000001101100000",
"111111111111101110111" when "000000000001110000000",
"111111111111110011011" when "000000000001110100000",
"111111111111110111101" when "000000000001111000000",
"111111111111111011111" when "000000000001111100000",
"000000000000000000000" when "000000000010000000000",
"000000000000000111110" when "000000000010001000000",
"000000000000001111000" when "000000000010010000000",
"000000000000010101111" when "000000000010011000000",
"000000000000011100100" when "000000000010100000000",
"000000000000100010110" when "000000000010101000000",
"000000000000101000110" when "000000000010110000000",
"000000000000101110011" when "000000000010111000000",
"000000000000110011111" when "000000000011000000000",
"000000000000111001000" when "000000000011001000000",
"000000000000111110001" when "000000000011010000000",
"000000000001000010111" when "000000000011011000000",
"000000000001000111101" when "000000000011100000000",
"000000000001001100000" when "000000000011101000000",
"000000000001010000011" when "000000000011110000000",
"000000000001010100101" when "000000000011111000000",
"000000000001011000101" when "000000000100000000000",
"000000000001100000011" when "000000000100010000000",
"000000000001100111110" when "000000000100100000000",
"000000000001101110101" when "000000000100110000000",
"000000000001110101010" when "000000000101000000000",
"000000000001111011100" when "000000000101010000000",
"000000000010000001011" when "000000000101100000000",
"000000000010000111001" when "000000000101110000000",
"000000000010001100100" when "000000000110000000000",
"000000000010010001110" when "000000000110010000000",
"000000000010010110110" when "000000000110100000000",
"000000000010011011101" when "000000000110110000000",
"000000000010100000010" when "000000000111000000000",
"000000000010100100110" when "000000000111010000000",
"000000000010101001001" when "000000000111100000000",
"000000000010101101011" when "000000000111110000000",
"000000000010110001011" when "000000001000000000000",
"000000000010111001001" when "000000001000100000000",
"000000000011000000100" when "000000001001000000000",
"000000000011000111011" when "000000001001100000000",
"000000000011001110000" when "000000001010000000000",
"000000000011010100010" when "000000001010100000000",
"000000000011011010001" when "000000001011000000000",
"000000000011011111111" when "000000001011100000000",
"000000000011100101010" when "000000001100000000000",
"000000000011101010100" when "000000001100100000000",
"000000000011101111100" when "000000001101000000000",
"000000000011110100011" when "000000001101100000000",
"000000000011111001000" when "000000001110000000000",
"000000000011111101100" when "000000001110100000000",
"000000000100000001111" when "000000001111000000000",
"000000000100000110000" when "000000001111100000000",
"000000000100001010001" when "000000010000000000000",
"000000000100010001111" when "000000010001000000000",
"000000000100011001001" when "000000010010000000000",
"000000000100100000001" when "000000010011000000000",
"000000000100100110101" when "000000010100000000000",
"000000000100101100111" when "000000010101000000000",
"000000000100110010111" when "000000010110000000000",
"000000000100111000100" when "000000010111000000000",
"000000000100111110000" when "000000011000000000000",
"000000000101000011010" when "000000011001000000000",
"000000000101001000010" when "000000011010000000000",
"000000000101001101001" when "000000011011000000000",
"000000000101010001110" when "000000011100000000000",
"000000000101010110010" when "000000011101000000000",
"000000000101011010101" when "000000011110000000000",
"000000000101011110110" when "000000011111000000000",
"000000000101100010111" when "000000100000000000000",


						"000000000000000000000" when others;
						
with valor select
	xlogmx 			<= 
"111111111111101110001" when "000000000000000100000",
"111111111111100001110" when "000000000000001000000",
"111111111111010111100" when "000000000000001100000",
"111111111111001110101" when "000000000000010000000",
"111111111111000110110" when "000000000000010100000",
"111111111110111111110" when "000000000000011000000",
"111111111110111001011" when "000000000000011100000",
"111111111110110011101" when "000000000000100000000",
"111111111110101110010" when "000000000000100100000",
"111111111110101001011" when "000000000000101000000",
"111111111110100101000" when "000000000000101100000",
"111111111110100000111" when "000000000000110000000",
"111111111110011101001" when "000000000000110100000",
"111111111110011001101" when "000000000000111000000",
"111111111110010110100" when "000000000000111100000",
"111111111110010011101" when "000000000001000000000",
"111111111110010000111" when "000000000001000100000",
"111111111110001110100" when "000000000001001000000",
"111111111110001100011" when "000000000001001100000",
"111111111110001010011" when "000000000001010000000",
"111111111110001000100" when "000000000001010100000",
"111111111110000111000" when "000000000001011000000",
"111111111110000101100" when "000000000001011100000",
"111111111110000100011" when "000000000001100000000",
"111111111110000011010" when "000000000001100100000",
"111111111110000010011" when "000000000001101000000",
"111111111110000001101" when "000000000001101100000",
"111111111110000001000" when "000000000001110000000",
"111111111110000000100" when "000000000001110100000",
"111111111110000000010" when "000000000001111000000",
"111111111110000000000" when "000000000001111100000",
"111111111110000000000" when "000000000010000000000",
"111111111110000000001" when "000000000010001000000",
"111111111110000000111" when "000000000010010000000",
"111111111110000010000" when "000000000010011000000",
"111111111110000011101" when "000000000010100000000",
"111111111110000101101" when "000000000010101000000",
"111111111110001000000" when "000000000010110000000",
"111111111110001010110" when "000000000010111000000",
"111111111110001101110" when "000000000011000000000",
"111111111110010001010" when "000000000011001000000",
"111111111110010100111" when "000000000011010000000",
"111111111110011001000" when "000000000011011000000",
"111111111110011101010" when "000000000011100000000",
"111111111110100001111" when "000000000011101000000",
"111111111110100110110" when "000000000011110000000",
"111111111110101100000" when "000000000011111000000",
"111111111110110001011" when "000000000100000000000",
"111111111110111101000" when "000000000100010000000",
"111111111111001001100" when "000000000100100000000",
"111111111111010110111" when "000000000100110000000",
"111111111111100101001" when "000000000101000000000",
"111111111111110100010" when "000000000101010000000",
"000000000000000100000" when "000000000101100000000",
"000000000000010100101" when "000000000101110000000",
"000000000000100101110" when "000000000110000000000",
"000000000000110111110" when "000000000110010000000",
"000000000001001010010" when "000000000110100000000",
"000000000001011101011" when "000000000110110000000",
"000000000001110001001" when "000000000111000000000",
"000000000010000101100" when "000000000111010000000",
"000000000010011010011" when "000000000111100000000",
"000000000010101111110" when "000000000111110000000",
"000000000011000101110" when "000000001000000000000",
"000000000011110011000" when "000000001000100000000",
"000000000100100010010" when "000000001001000000000",
"000000000101010011010" when "000000001001100000000",
"000000000110000110000" when "000000001010000000000",
"000000000110111010010" when "000000001010100000000",
"000000000111110000001" when "000000001011000000000",
"000000001000100111011" when "000000001011100000000",
"000000001001100000000" when "000000001100000000000",
"000000001010011010000" when "000000001100100000000",
"000000001011010101010" when "000000001101000000000",
"000000001100010001110" when "000000001101100000000",
"000000001101001111100" when "000000001110000000000",
"000000001110001110010" when "000000001110100000000",
"000000001111001110010" when "000000001111000000000",
"000000010000001111010" when "000000001111100000000",
"000000010001010001010" when "000000010000000000000",
"000000010011011000011" when "000000010001000000000",
"000000010101100011001" when "000000010010000000000",
"000000010111110001100" when "000000010011000000000",
"000000011010000011010" when "000000010100000000000",
"000000011100011000001" when "000000010101000000000",
"000000011110110000001" when "000000010110000000000",
"000000100001001011001" when "000000010111000000000",
"000000100011101000110" when "000000011000000000000",
"000000100110001001001" when "000000011001000000000",
"000000101000101100000" when "000000011010000000000",
"000000101011010001011" when "000000011011000000000",
"000000101101111001001" when "000000011100000000000",
"000000110000100011001" when "000000011101000000000",
"000000110011001111011" when "000000011110000000000",
"000000110101111101110" when "000000011111000000000",
"000000111000101110010" when "000000100000000000000",
						"000000000000000000000" when others;


end Behavioral;


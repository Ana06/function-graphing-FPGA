----------------------------------------------------------------------------------
-- Company: Nameless2
-- Engineer: Ana María Martínez Gómez, Aitor Alonso Lorenzo, Víctor Adolfo Gallego Alcalá
-- 
-- Create Date:    13:18:25 02/19/2014 
-- Design Name: 
-- Module Name:    trigo - Behavioral 
-- Project Name: Representación gráfica de funciones	
-- Target Devices: 
-- Tool versions: 
-- Description: 
--
-- Dependencies: 
--
-- Revision: 
-- Revision 0.01 - File Created
-- Additional Comments: 
--
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity trigo is
    Port ( valor : in  STD_LOGIC_VECTOR (20 downto 0);
           sen : out  STD_LOGIC_VECTOR (20 downto 0);
           cos : out  STD_LOGIC_VECTOR (20 downto 0));
end trigo;

architecture Behavioral of trigo is

begin

with valor select
	sen 	<= 		"000000000000000000000" when "111111100000000000000",
"111111111111111111111" when "111111100010000000000",
"000000000000000000000" when "111111100100000000000",
"000000000000000000000" when "111111100110000000000",
"000000000000000000000" when "111111101000000000000",
"111111111111111111111" when "111111101010000000000",
"000000000000000000000" when "111111101100000000000",
"111111111111111111111" when "111111101110000000000",
"000000000000000000000" when "111111110000000000000",
"000000000010000000000" when "111111110001000000000",
"111111111111111111111" when "111111110010000000000",
"111111111110000000000" when "111111110011000000000",
"000000000000000000000" when "111111110100000000000",
"000000000010000000000" when "111111110101000000000",
"111111111111111111111" when "111111110110000000000",
"111111111110000000000" when "111111110111000000000",
"000000000000000000000" when "111111111000000000000",
"000000000001011010100" when "111111111000100000000",
"000000000010000000000" when "111111111001000000000",
"000000000001011010100" when "111111111001100000000",
"111111111111111111111" when "111111111010000000000",
"111111111110100101011" when "111111111010100000000",
"111111111110000000000" when "111111111011000000000",
"111111111110100101011" when "111111111011100000000",
"000000000000000000000" when "111111111100000000000",
"000000000000110000111" when "111111111100010000000",
"000000000001011010100" when "111111111100100000000",
"000000000001110110010" when "111111111100110000000",
"000000000010000000000" when "111111111101000000000",
"000000000001110110010" when "111111111101010000000",
"000000000001011010100" when "111111111101100000000",
"000000000000110000111" when "111111111101110000000",
"111111111111111111111" when "111111111110000000000",
"111111111111100111000" when "111111111110001000000",
"111111111111001111000" when "111111111110010000000",
"111111111110111000111" when "111111111110011000000",
"111111111110100101011" when "111111111110100000000",
"111111111110010101100" when "111111111110101000000",
"111111111110001001101" when "111111111110110000000",
"111111111110000010011" when "111111111110111000000",
"111111111110000000000" when "111111111111000000000",
"111111111110000010011" when "111111111111001000000",
"111111111110001001101" when "111111111111010000000",
"111111111110010101100" when "111111111111011000000",
"111111111110100101011" when "111111111111100000000",
"111111111110111000111" when "111111111111101000000",
"111111111111001111000" when "111111111111110000000",
"111111111111100111000" when "111111111111111000000",
"000000000000000000000" when "000000000000000000000",
"000000000000001100100" when "000000000000000100000",
"000000000000011000111" when "000000000000001000000",
"000000000000100101001" when "000000000000001100000",
"000000000000110000111" when "000000000000010000000",
"000000000000111100010" when "000000000000010100000",
"000000000001000111000" when "000000000000011000000",
"000000000001010001001" when "000000000000011100000",
"000000000001011010100" when "000000000000100000000",
"000000000001100010111" when "000000000000100100000",
"000000000001101010011" when "000000000000101000000",
"000000000001110000111" when "000000000000101100000",
"000000000001110110010" when "000000000000110000000",
"000000000001111010011" when "000000000000110100000",
"000000000001111101100" when "000000000000111000000",
"000000000001111111011" when "000000000000111100000",
"000000000010000000000" when "000000000001000000000",
"000000000001111111011" when "000000000001000100000",
"000000000001111101100" when "000000000001001000000",
"000000000001111010011" when "000000000001001100000",
"000000000001110110010" when "000000000001010000000",
"000000000001110000111" when "000000000001010100000",
"000000000001101010011" when "000000000001011000000",
"000000000001100010111" when "000000000001011100000",
"000000000001011010100" when "000000000001100000000",
"000000000001010001001" when "000000000001100100000",
"000000000001000111000" when "000000000001101000000",
"000000000000111100010" when "000000000001101100000",
"000000000000110000111" when "000000000001110000000",
"000000000000100101001" when "000000000001110100000",
"000000000000011000111" when "000000000001111000000",
"000000000000001100100" when "000000000001111100000",
"000000000000000000000" when "000000000010000000000",
"111111111111100111000" when "000000000010001000000",
"111111111111001111000" when "000000000010010000000",
"111111111110111000111" when "000000000010011000000",
"111111111110100101011" when "000000000010100000000",
"111111111110010101100" when "000000000010101000000",
"111111111110001001101" when "000000000010110000000",
"111111111110000010011" when "000000000010111000000",
"111111111110000000000" when "000000000011000000000",
"111111111110000010011" when "000000000011001000000",
"111111111110001001101" when "000000000011010000000",
"111111111110010101100" when "000000000011011000000",
"111111111110100101011" when "000000000011100000000",
"111111111110111000111" when "000000000011101000000",
"111111111111001111000" when "000000000011110000000",
"111111111111100111000" when "000000000011111000000",
"111111111111111111111" when "000000000100000000000",
"000000000000110000111" when "000000000100010000000",
"000000000001011010100" when "000000000100100000000",
"000000000001110110010" when "000000000100110000000",
"000000000010000000000" when "000000000101000000000",
"000000000001110110010" when "000000000101010000000",
"000000000001011010100" when "000000000101100000000",
"000000000000110000111" when "000000000101110000000",
"000000000000000000000" when "000000000110000000000",
"111111111111001111000" when "000000000110010000000",
"111111111110100101011" when "000000000110100000000",
"111111111110001001101" when "000000000110110000000",
"111111111110000000000" when "000000000111000000000",
"111111111110001001101" when "000000000111010000000",
"111111111110100101011" when "000000000111100000000",
"111111111111001111000" when "000000000111110000000",
"111111111111111111111" when "000000001000000000000",
"000000000001011010100" when "000000001000100000000",
"000000000010000000000" when "000000001001000000000",
"000000000001011010100" when "000000001001100000000",
"000000000000000000000" when "000000001010000000000",
"111111111110100101011" when "000000001010100000000",
"111111111110000000000" when "000000001011000000000",
"111111111110100101011" when "000000001011100000000",
"111111111111111111111" when "000000001100000000000",
"000000000001011010100" when "000000001100100000000",
"000000000010000000000" when "000000001101000000000",
"000000000001011010100" when "000000001101100000000",
"000000000000000000000" when "000000001110000000000",
"111111111110100101011" when "000000001110100000000",
"111111111110000000000" when "000000001111000000000",
"111111111110100101011" when "000000001111100000000",
"111111111111111111111" when "000000010000000000000",
"000000000010000000000" when "000000010001000000000",
"000000000000000000000" when "000000010010000000000",
"111111111110000000000" when "000000010011000000000",
"111111111111111111111" when "000000010100000000000",
"000000000010000000000" when "000000010101000000000",
"000000000000000000000" when "000000010110000000000",
"111111111110000000000" when "000000010111000000000",
"111111111111111111111" when "000000011000000000000",
"000000000010000000000" when "000000011001000000000",
"111111111111111111111" when "000000011010000000000",
"111111111110000000000" when "000000011011000000000",
"111111111111111111111" when "000000011100000000000",
"000000000010000000000" when "000000011101000000000",
"000000000000000000000" when "000000011110000000000",
"111111111110000000000" when "000000011111000000000",
"111111111111111111111" when "000000100000000000000",


						"000000000000000000000" when others;
						
with valor select
	cos		 	<= "000000000010000000000" when "111111100000000000000",
"111111111110000000000" when "111111100010000000000",
"000000000010000000000" when "111111100100000000000",
"111111111110000000000" when "111111100110000000000",
"000000000010000000000" when "111111101000000000000",
"111111111110000000000" when "111111101010000000000",
"000000000010000000000" when "111111101100000000000",
"111111111110000000000" when "111111101110000000000",
"000000000010000000000" when "111111110000000000000",
"111111111111111111111" when "111111110001000000000",
"111111111110000000000" when "111111110010000000000",
"111111111111111111111" when "111111110011000000000",
"000000000010000000000" when "111111110100000000000",
"111111111111111111111" when "111111110101000000000",
"111111111110000000000" when "111111110110000000000",
"000000000000000000000" when "111111110111000000000",
"000000000010000000000" when "111111111000000000000",
"000000000001011010100" when "111111111000100000000",
"111111111111111111111" when "111111111001000000000",
"111111111110100101011" when "111111111001100000000",
"111111111110000000000" when "111111111010000000000",
"111111111110100101011" when "111111111010100000000",
"000000000000000000000" when "111111111011000000000",
"000000000001011010100" when "111111111011100000000",
"000000000010000000000" when "111111111100000000000",
"000000000001110110010" when "111111111100010000000",
"000000000001011010100" when "111111111100100000000",
"000000000000110000111" when "111111111100110000000",
"111111111111111111111" when "111111111101000000000",
"111111111111001111000" when "111111111101010000000",
"111111111110100101011" when "111111111101100000000",
"111111111110001001101" when "111111111101110000000",
"111111111110000000000" when "111111111110000000000",
"111111111110000010011" when "111111111110001000000",
"111111111110001001101" when "111111111110010000000",
"111111111110010101100" when "111111111110011000000",
"111111111110100101011" when "111111111110100000000",
"111111111110111000111" when "111111111110101000000",
"111111111111001111000" when "111111111110110000000",
"111111111111100111000" when "111111111110111000000",
"000000000000000000000" when "111111111111000000000",
"000000000000011000111" when "111111111111001000000",
"000000000000110000111" when "111111111111010000000",
"000000000001000111000" when "111111111111011000000",
"000000000001011010100" when "111111111111100000000",
"000000000001101010011" when "111111111111101000000",
"000000000001110110010" when "111111111111110000000",
"000000000001111101100" when "111111111111111000000",
"000000000010000000000" when "000000000000000000000",
"000000000001111111011" when "000000000000000100000",
"000000000001111101100" when "000000000000001000000",
"000000000001111010011" when "000000000000001100000",
"000000000001110110010" when "000000000000010000000",
"000000000001110000111" when "000000000000010100000",
"000000000001101010011" when "000000000000011000000",
"000000000001100010111" when "000000000000011100000",
"000000000001011010100" when "000000000000100000000",
"000000000001010001001" when "000000000000100100000",
"000000000001000111000" when "000000000000101000000",
"000000000000111100010" when "000000000000101100000",
"000000000000110000111" when "000000000000110000000",
"000000000000100101001" when "000000000000110100000",
"000000000000011000111" when "000000000000111000000",
"000000000000001100100" when "000000000000111100000",
"000000000000000000000" when "000000000001000000000",
"111111111111110011011" when "000000000001000100000",
"111111111111100111000" when "000000000001001000000",
"111111111111011010110" when "000000000001001100000",
"111111111111001111000" when "000000000001010000000",
"111111111111000011101" when "000000000001010100000",
"111111111110111000111" when "000000000001011000000",
"111111111110101110110" when "000000000001011100000",
"111111111110100101011" when "000000000001100000000",
"111111111110011101000" when "000000000001100100000",
"111111111110010101100" when "000000000001101000000",
"111111111110001111000" when "000000000001101100000",
"111111111110001001101" when "000000000001110000000",
"111111111110000101100" when "000000000001110100000",
"111111111110000010011" when "000000000001111000000",
"111111111110000000100" when "000000000001111100000",
"111111111110000000000" when "000000000010000000000",
"111111111110000010011" when "000000000010001000000",
"111111111110001001101" when "000000000010010000000",
"111111111110010101100" when "000000000010011000000",
"111111111110100101011" when "000000000010100000000",
"111111111110111000111" when "000000000010101000000",
"111111111111001111000" when "000000000010110000000",
"111111111111100111000" when "000000000010111000000",
"111111111111111111111" when "000000000011000000000",
"000000000000011000111" when "000000000011001000000",
"000000000000110000111" when "000000000011010000000",
"000000000001000111000" when "000000000011011000000",
"000000000001011010100" when "000000000011100000000",
"000000000001101010011" when "000000000011101000000",
"000000000001110110010" when "000000000011110000000",
"000000000001111101100" when "000000000011111000000",
"000000000010000000000" when "000000000100000000000",
"000000000001110110010" when "000000000100010000000",
"000000000001011010100" when "000000000100100000000",
"000000000000110000111" when "000000000100110000000",
"000000000000000000000" when "000000000101000000000",
"111111111111001111000" when "000000000101010000000",
"111111111110100101011" when "000000000101100000000",
"111111111110001001101" when "000000000101110000000",
"111111111110000000000" when "000000000110000000000",
"111111111110001001101" when "000000000110010000000",
"111111111110100101011" when "000000000110100000000",
"111111111111001111000" when "000000000110110000000",
"111111111111111111111" when "000000000111000000000",
"000000000000110000111" when "000000000111010000000",
"000000000001011010100" when "000000000111100000000",
"000000000001110110010" when "000000000111110000000",
"000000000010000000000" when "000000001000000000000",
"000000000001011010100" when "000000001000100000000",
"000000000000000000000" when "000000001001000000000",
"111111111110100101011" when "000000001001100000000",
"111111111110000000000" when "000000001010000000000",
"111111111110100101011" when "000000001010100000000",
"111111111111111111111" when "000000001011000000000",
"000000000001011010100" when "000000001011100000000",
"000000000010000000000" when "000000001100000000000",
"000000000001011010100" when "000000001100100000000",
"111111111111111111111" when "000000001101000000000",
"111111111110100101011" when "000000001101100000000",
"111111111110000000000" when "000000001110000000000",
"111111111110100101011" when "000000001110100000000",
"111111111111111111111" when "000000001111000000000",
"000000000001011010100" when "000000001111100000000",
"000000000010000000000" when "000000010000000000000",
"111111111111111111111" when "000000010001000000000",
"111111111110000000000" when "000000010010000000000",
"111111111111111111111" when "000000010011000000000",
"000000000010000000000" when "000000010100000000000",
"111111111111111111111" when "000000010101000000000",
"111111111110000000000" when "000000010110000000000",
"111111111111111111111" when "000000010111000000000",
"000000000010000000000" when "000000011000000000000",
"111111111111111111111" when "000000011001000000000",
"111111111110000000000" when "000000011010000000000",
"111111111111111111111" when "000000011011000000000",
"000000000010000000000" when "000000011100000000000",
"111111111111111111111" when "000000011101000000000",
"111111111110000000000" when "000000011110000000000",
"111111111111111111111" when "000000011111000000000",
"000000000010000000000" when "000000100000000000000",


						"000000000000000000000" when others;


end Behavioral;

